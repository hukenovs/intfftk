-------------------------------------------------------------------------------
--
-- Title       : iobuf_two_rw
-- Design      : fpfftk
-- Author      : Kapitanov
-- Company     :
--
-------------------------------------------------------------------------------
--
-- Description : version 1.0
--
-------------------------------------------------------------------------------
--
--	Version 1.0  12.02.2016
--        Description: Convert data from interleave-2 mode to bit-reverse.
--                        Common clock. Input data enable strobe CAN be wrapped! 
--                        
--        Example 1 (Mode BITREV = FALSE): Interleave-2 to Half-part data.		
--
--        Data in:
--            DIx: ...0246...
--            DIx: ...1357...
--
--        Data out: (two parts of data)
--            DOx: .......0123...
--            DOx: .......4567...
--
--        Example 2 (Mode BITREV = TRUE): Half-part data to Interleave-2.		
--
--        Data in:
--            DIx: ...0123...
--            DIx: ...4567...
--
--        Data out: (interleave-2)
--            DOx: .......0246...
--            DOx: .......1357...
--
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
--
--	GNU GENERAL PUBLIC LICENSE
--  Version 3, 29 June 2007
--
--	Copyright (c) 2018 Kapitanov Alexander
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--  THERE IS NO WARRANTY FOR THE PROGRAM, TO THE EXTENT PERMITTED BY
--  APPLICABLE LAW. EXCEPT WHEN OTHERWISE STATED IN WRITING THE COPYRIGHT 
--  HOLDERS AND/OR OTHER PARTIES PROVIDE THE PROGRAM "AS IS" WITHOUT WARRANTY 
--  OF ANY KIND, EITHER EXPRESSED OR IMPLIED, INCLUDING, BUT NOT LIMITED TO, 
--  THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR 
--  PURPOSE.  THE ENTIRE RISK AS TO THE QUALITY AND PERFORMANCE OF THE PROGRAM 
--  IS WITH YOU.  SHOULD THE PROGRAM PROVE DEFECTIVE, YOU ASSUME THE COST OF 
--  ALL NECESSARY SERVICING, REPAIR OR CORRECTION. 
-- 
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity iobuf_two_rw is
	generic (
		TD			: time:=0.1ns;   --! Simulation time
		BITREV		: boolean:=FALSE;--! Bit-reverse mode (FALSE - int2-to-half, TRUE - half-to-int2)
		DATA		: integer:= 32;  --! Data Width
	    ADDR		: integer:= 10   --! Address depth
		);
	port (
	    rst			: in  std_logic; --! Common reset (high)
		clk			: in  std_logic; --! Common clock	    

	    dt_int0		: in  std_logic_vector(DATA-1 downto 0);    
	    dt_int1		: in  std_logic_vector(DATA-1 downto 0);    
	    dt_en01		: in  std_logic;
		
	    dt_rev0		: out std_logic_vector(DATA-1 downto 0);
	    dt_rev1		: out std_logic_vector(DATA-1 downto 0);
		dt_vl01		: out std_logic
	);
end iobuf_two_rw;
 
architecture iobuf_two_rw of iobuf_two_rw is

---------------- Calculate Index Counter ----------------
type add_type is array(0 to ADDR-1) of std_logic_vector(ADDR-2 downto 0);
type inc_type is array(0 to ADDR-1) of std_logic_vector(ADDR-2 downto 0);
type msb_type is array(0 to ADDR-1) of integer;

function adr_msb return msb_type is
	variable tmp_ret : msb_type;
begin
	tmp_ret(0) := ADDR-1;
	xL: for ii in 1 to ADDR-1 loop
		tmp_ret(ii) := ii-1;
	end loop;
	return tmp_ret;
end function;

function adr_shift return inc_type is
	variable tmp_arr : std_logic_vector(ADDR-1 downto 0);
	variable tmp_ret : inc_type;
begin
	xL: for ii in 0 to ADDR-1 loop
		tmp_arr := ((ADDR-1-ii) => '1', others => '0');
		tmp_ret(ii) := tmp_arr(ADDR-2 downto 0);
	end loop;

	return tmp_ret;
end function;

function adr_increment return add_type is
	variable tmp_arr : std_logic_vector(ADDR-1 downto 0);
	variable tmp_ret : add_type;
begin
	tmp_ret(0) := (0 => '1', others => '0');
	xL: for ii in 1 to ADDR-1 loop
		tmp_arr :=  ((ADDR-ii) => '1', others => '0');
		tmp_ret(ii) := tmp_arr(ADDR-2 downto 0);
	end loop;
	return tmp_ret;
end function;

constant INC_MSB 		: msb_type:=adr_msb; 
constant INC_DEL 		: inc_type:=adr_shift; 
constant INC_ADD 		: add_type:=adr_increment;
 
---------------- Write / Read pointers ----------------
signal WR_MSB			: integer range 0 to ADDR-1;
signal WR_DEL			: std_logic_vector(ADDR-2 downto 0);
signal WR_ADD			: std_logic_vector(ADDR-2 downto 0);

signal RD_MSB			: integer range 0 to ADDR-1;
signal RD_DEL			: std_logic_vector(ADDR-2 downto 0);
signal RD_ADD			: std_logic_vector(ADDR-2 downto 0);

signal RD_INZ			: std_logic_vector(ADDR-2 downto 0);
signal WR_INZ			: std_logic_vector(ADDR-2 downto 0);


signal dt_ena			: std_logic;

---------------- RAM signals ----------------
signal ram_dia			: std_logic_vector(DATA-1 downto 0);
signal ram_dib			: std_logic_vector(DATA-1 downto 0);
	
signal ram0_dia			: std_logic_vector(DATA-1 downto 0);
signal ram0_dib			: std_logic_vector(DATA-1 downto 0);
signal ram1_dia			: std_logic_vector(DATA-1 downto 0);
signal ram1_dib			: std_logic_vector(DATA-1 downto 0);

signal ram0_doa			: std_logic_vector(DATA-1 downto 0);
signal ram0_dob			: std_logic_vector(DATA-1 downto 0);
signal ram1_doa			: std_logic_vector(DATA-1 downto 0);
signal ram1_dob			: std_logic_vector(DATA-1 downto 0);

---------------- Calculate Bit / Index Position -----------------
signal sw_inc			: std_logic;
signal sw_ena			: std_logic;

signal cnt_even			: std_logic_vector(ADDR-1 downto 0);
signal cnt_odd			: std_logic_vector(ADDR-1 downto 0);
signal sw_ptr			: std_logic_vector(ADDR-1 downto 0);



signal in_cnt			: integer range 0 to ADDR-1;
signal sw_cnt			: std_logic_vector(ADDR-1 downto 0);
signal sw_adr			: std_logic_vector(ADDR-1 downto 0);

signal cnt_wr0			: std_logic_vector(ADDR-2 downto 0);
signal cnt_wr1			: std_logic_vector(ADDR-2 downto 0);
signal cnt_rd0			: std_logic_vector(ADDR-2 downto 0);
signal cnt_rd1			: std_logic_vector(ADDR-2 downto 0);

signal adr_wr0			: std_logic_vector(ADDR-2 downto 0);
signal adr_wr1			: std_logic_vector(ADDR-2 downto 0);
signal adr_rd0			: std_logic_vector(ADDR-2 downto 0);
signal adr_rd1			: std_logic_vector(ADDR-2 downto 0);

signal ram0_wr0			: std_logic;
signal ram0_wr1			: std_logic;
signal ram1_wr0			: std_logic;
signal ram1_wr1			: std_logic;

signal ram0_we0			: std_logic;
signal ram0_we1			: std_logic;
signal ram1_we0			: std_logic;
signal ram1_we1			: std_logic;

signal ram0_rd0			: std_logic;
signal ram0_rd1			: std_logic;
signal ram1_rd0			: std_logic;
signal ram1_rd1			: std_logic;

signal cnt_ptr			: std_logic_vector(ADDR-1 downto 0);
signal cnt_ena			: std_logic;

begin

---------------- Write Increment ---------------- 
pr_del: process(clk) is
begin
	if rising_edge(clk) then
		if (rst = '1') then
			sw_cnt <= (0 => '1', others => '0') after td;
			sw_adr <= (others => '0') after td;

			in_cnt <= 1 after td;
			WR_MSB <= INC_MSB(0) after td;
			WR_DEL <= INC_DEL(0) after td;
			WR_ADD <= INC_ADD(0) after td;
		else
			if (dt_en01 = '1') then				
				sw_adr <= sw_adr + '1' after td;
				---- Counter for WR0 / WR1 ----
				if (sw_cnt(sw_cnt'left) = '1') then
					sw_cnt <= (0 => '1', others => '0') after td;
				else
					sw_cnt <= sw_cnt + '1' after td;
				end if;					

				---- Counter for Arrays ----
				if (sw_cnt(sw_cnt'left) = '1') then	
					if (in_cnt = (ADDR-1)) then
						in_cnt <= 0 after td;
					else
						in_cnt <= in_cnt + 1 after td;
					end if;
					WR_MSB <= INC_MSB(in_cnt) after td;
					WR_DEL <= INC_DEL(in_cnt) after td;
					WR_ADD <= INC_ADD(in_cnt) after td;
				end if;						
			end if;	
			sw_inc <= sw_cnt(sw_cnt'left) after td;
		end if;
	end if;
end process;

WR_INZ <= WR_ADD after td when rising_edge(clk);

---------------- Write Counters ---------------- 
pr_wr: process(clk) is
begin
	if rising_edge(clk) then
		dt_ena <= dt_en01 after td;
		
		if (rst = '1') then
			ram0_wr0 <= '0' after td;
			ram0_wr1 <= '0' after td;
			ram1_wr0 <= '0' after td;
			ram1_wr1 <= '0' after td;
			
			cnt_wr0 <= (others => '0') after td;
			cnt_wr1 <= WR_DEL after td;

			cnt_ptr <= (0 => '1', others => '0') after td;
			cnt_ena	<= '0' after td;
		else
			---- Write enable ----
			if (dt_en01 = '1') then
				if (cnt_ptr(WR_MSB) = '1') then
					cnt_ptr <= (0 => '1', others => '0') after td;
					cnt_ena <= '1' after td;
				else
					cnt_ptr <= cnt_ptr + '1' after td;
					cnt_ena <= '0' after td;
				end if;
			end if;	
			
			---- Find increment mux ----
			if (dt_en01 = '1') then
				ram0_wr0 <= not sw_adr(WR_MSB) after td;
				ram0_wr1 <= not (WR_ADD(0) or sw_adr(WR_MSB)) after td;
				ram1_wr0 <= WR_ADD(0) or sw_adr(WR_MSB) after td;
				ram1_wr1 <= not WR_ADD(0) and sw_adr(WR_MSB) after td;
			end if;			

			---- Find adress counter ----
			if (dt_ena = '1') then		
				if (sw_inc = '1') then
					cnt_wr0 <= (others => '0') after td;
					cnt_wr1 <= WR_DEL after td;
				else
					---- Write Counter ----
					if (cnt_ena = '1' and ram0_wr1 = '0') then
						cnt_wr0 <= cnt_wr0 + WR_INZ + 1 after td;
						cnt_wr1 <= cnt_wr1 + WR_INZ + 1 after td;
					else
						cnt_wr0 <= cnt_wr0 + WR_INZ after td;
						cnt_wr1 <= cnt_wr1 + WR_INZ after td;
					end if;						
					
				end if;	
			end if;
		end if;
	end if;
end process;

---- RAM 0/1 mapping ----
pr_din: process(clk) is
begin
	if rising_edge(clk) then
		---- Input data delays ----
		ram_dia <= dt_int0 after td;
		ram_dib <= dt_int1 after td;
		---- Mux input data ----
		if (ram0_wr0 = '1') then
			ram0_dia <= ram_dia after td;
            ram0_dib <= ram_dib after td;
		end if;
		if (ram1_wr0 = '1') then
			ram1_dia <= ram_dib after td;
            ram1_dib <= ram_dia after td;
		end if;
		---- Write enable to RAMBs ----
		ram0_we0 <= ram0_wr0 after td;
		ram0_we1 <= ram0_wr1 after td;
		ram1_we0 <= ram1_wr0 after td;
		ram1_we1 <= ram1_wr1 after td;
		---- Address R/W RAMBs ----
		adr_wr0 <= cnt_wr0 after td;
		adr_wr1 <= cnt_wr1 after td;
		adr_rd0 <= cnt_rd0 after td;
		adr_rd1 <= cnt_rd1 after td;
	end if;
end process;

-- xTDP_RAM0: entity work.ramb_tdp_rw
	-- generic map (
	    -- DATA    => DATA,
	    -- ADDR    => ADDR-1
		-- )
	-- port map (
		-- clk     => clk,
		-- -- Port A --
	    -- a_wr    => ram0_wr0,
	    -- a_rd    => ram_rd,
		-- a_adr   => adr_wr0,
	    -- a_din   => ram0_dia, 
	    -- a_dout  => ram_doa,
	    -- -- Port B --
	    -- b_wr    => ram0_wr1,
	    -- b_rd    => ram_rd,
		-- b_adr   => adr_wr1,
	    -- b_din   => ram0_dib, 
	    -- b_dout  => ram_dob
	-- );

-- xTDP_RAM1: entity work.ramb_tdp_rw
	-- generic map (
	    -- DATA    => DATA,
	    -- ADDR    => ADDR-1
		-- )
	-- port map (
		-- clk     => clk,
		-- -- Port A --
	    -- a_wr    => ram1_wr0,
	    -- a_rd    => ram_rd,
		-- a_adr   => adr_wr0,
	    -- a_din   => ram1_dia, 
	    -- a_dout  => ram_doa,
	    -- -- Port B --
	    -- b_wr    => ram1_wr1,
	    -- b_rd    => ram_rd,
		-- b_adr   => adr_wr1,
	    -- b_din   => ram1_dib, 
	    -- b_dout  => ram_dob
	-- );
	
	
end iobuf_two_rw;